module light_up();
    
endmodule